library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Ensamblado is
    Port ( clr,clr : in  STD_LOGIC;
           datos : out  STD_LOGIC_VECTOR (7 downto 0));
end Ensamblado;

architecture Behavioral of Ensamblado is

begin


end Behavioral;

