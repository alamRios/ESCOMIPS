library IEEE;
use IEEE.STD_LOGIC_1164.all;

package ESCOMIPS_PAK is
end ESCOMIPS_PAK;

package body ESCOMIPS_PAK is
 
end ESCOMIPS_PAK;
